// $Id: $
// File name:   sensor_s.sv
// Created:     1/18/2023
// Author:      Wen-Bo Hung
// Lab Section: 337-04
// Version:     1.0  Initial Design Entry
// Description: Structural Style Sensor Error Detector.
